// 
//  Copyright 2022 Sergey Khabarov, sergeykhbr@gmail.com
// 
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
// 

`timescale 1ns/10ps

module pcie_io_rx_engine #(
    parameter int C_DATA_WIDTH = 64,
    parameter int KEEP_WIDTH = (C_DATA_WIDTH / 8)
)
(
    input logic i_nrst,
    input logic i_clk,                                      // System bus clock
    // 
    input logic [C_DATA_WIDTH-1:0] i_m_axis_rx_tdata,
    input logic [KEEP_WIDTH-1:0] i_m_axis_rx_tkeep,
    input logic i_m_axis_rx_tlast,
    input logic i_m_axis_rx_tvalid,
    output logic o_m_axis_rx_tready,
    input logic [8:0] i_m_axis_rx_tuser,
    // 
    output logic o_req_compl,
    output logic o_req_compl_wd,                            // req completion without data (IO WR32 request)
    input logic i_compl_done,
    // 
    output logic [2:0] o_req_tc,                            // Memory Read TC
    output logic o_req_td,                                  // Memory Read TD
    output logic o_req_ep,                                  // Memory Read EP
    output logic [1:0] o_req_attr,                          // Memory Read Attribute
    output logic [9:0] o_req_len,                           // Memory Read Length (1DW)
    output logic [15:0] o_req_rid,                          // Memory Read Requestor ID
    output logic [7:0] o_req_tag,                           // Memory Read Tag
    output logic [7:0] o_req_be,                            // Memory Read Byte Enables
    output logic [12:0] o_req_addr,                         // Memory Read Address
    // 
    input logic i_req_mem_ready,                            // Ready to accept next memory request
    output logic o_req_mem_valid,                           // Request data is valid to accept
    output logic o_req_mem_64,                              // 0=32-bits; 1=64-bits
    output logic o_req_mem_write,                           // 0=read; 1=write operation
    output logic [9:0] o_req_mem_bytes,                     // 0=1024 B; 4=DWORD; 8=QWORD; ...
    output logic [12:0] o_req_mem_addr,                     // Address to read/write
    output logic [7:0] o_req_mem_strob,                     // Byte enabling write strob
    output logic [63:0] o_req_mem_data,                     // Data to write
    output logic o_req_mem_last,                            // Last data payload in a sequence
    input logic i_resp_mem_valid                            // Read/Write data is valid. All write transaction with valid response.
);


localparam bit [6:0] PIO_RX_MEM_RD32_FMT_TYPE = 7'h00;
localparam bit [6:0] PIO_RX_MEM_WR32_FMT_TYPE = 7'h40;
localparam bit [6:0] PIO_RX_MEM_RD64_FMT_TYPE = 7'h20;
localparam bit [6:0] PIO_RX_MEM_WR64_FMT_TYPE = 7'h60;
localparam bit [6:0] PIO_RX_IO_RD32_FMT_TYPE = 7'h02;
localparam bit [6:0] PIO_RX_IO_WR32_FMT_TYPE = 7'h42;

localparam bit [7:0] PIO_RX_RST_STATE = 8'h00;
localparam bit [7:0] PIO_RX_MEM_RD32_DW1DW2 = 8'h01;
localparam bit [7:0] PIO_RX_MEM_WR32_DW1DW2 = 8'h02;
localparam bit [7:0] PIO_RX_MEM_RD64_DW1DW2 = 8'h04;
localparam bit [7:0] PIO_RX_MEM_WR64_DW1DW2 = 8'h08;
localparam bit [7:0] PIO_RX_MEM_WR64_DW3 = 8'h10;
localparam bit [7:0] PIO_RX_IO_WR_DW1DW2 = 8'h20;
localparam bit [7:0] PIO_RX_WAIT_DMA_RESP = 8'h40;
localparam bit [7:0] PIO_RX_WAIT_TX_COMPLETION = 8'h80;
// TLP Response Types:
localparam bit [1:0] TLP_NON_POSTED = 2'd0;                 // No response at all
localparam bit [1:0] TLP_POSTED = 2'd3;                     // Response with data payload
localparam bit [1:0] TLP_COMPLETION = 2'd1;                 // Response without payload

typedef struct {
    logic m_axis_rx_tready;
    logic req_valid;
    logic [2:0] req_tc;
    logic req_td;
    logic req_ep;
    logic [1:0] req_attr;
    logic [9:0] req_len;
    logic [15:0] req_rid;
    logic [7:0] req_tag;
    logic [7:0] req_be;
    logic [12:0] req_addr;
    logic [10:0] wr_addr;
    logic [7:0] wr_be;
    logic wr_en;
    logic [63:0] wr_data;
    logic [7:0] state;
    logic [7:0] tlp_type;
    logic [1:0] tlp_resp;
} pcie_io_rx_engine_registers;

const pcie_io_rx_engine_registers pcie_io_rx_engine_r_reset = '{
    1'b0,                               // m_axis_rx_tready
    1'b0,                               // req_valid
    3'd0,                               // req_tc
    1'b0,                               // req_td
    1'b0,                               // req_ep
    2'd0,                               // req_attr
    10'd0,                              // req_len
    16'd0,                              // req_rid
    8'd0,                               // req_tag
    8'd0,                               // req_be
    13'd0,                              // req_addr
    11'd0,                              // wr_addr
    8'd0,                               // wr_be
    1'b0,                               // wr_en
    64'd0,                              // wr_data
    PIO_RX_RST_STATE,                   // state
    8'd0,                               // tlp_type
    TLP_NON_POSTED                      // tlp_resp
};
pcie_io_rx_engine_registers r;
pcie_io_rx_engine_registers rin;


always_comb
begin: comb_proc
    pcie_io_rx_engine_registers v;
    logic [1:0] vb_region_select;

    v = r;
    vb_region_select = '0;


    if (i_m_axis_rx_tuser[8: 2] == 7'h01) begin             // Select Mem32 region
        vb_region_select = 2'h1;
    end else if (i_m_axis_rx_tuser[8: 2] == 7'h02) begin    // Select Mem64 region
        vb_region_select = 2'h2;
    end else if (i_m_axis_rx_tuser[8: 2] == 7'h40) begin    // Select EROM region
        vb_region_select = 2'h3;
    end

    v.wr_en = 1'b0;

    case (r.state)
    PIO_RX_RST_STATE: begin
        v.m_axis_rx_tready = 1'b1;
        v.tlp_resp = 2'd0;

        if (i_m_axis_rx_tvalid == 1'b1) begin
            v.tlp_type = i_m_axis_rx_tdata[31: 24];
            v.req_len = i_m_axis_rx_tdata[9: 0];

            case (i_m_axis_rx_tdata[30: 24])
            PIO_RX_MEM_RD32_FMT_TYPE: begin
                if (i_m_axis_rx_tdata[9: 0] == 10'd1) begin
                    v.req_tc = i_m_axis_rx_tdata[22: 20];
                    v.req_td = i_m_axis_rx_tdata[15];
                    v.req_ep = i_m_axis_rx_tdata[14];
                    v.req_attr = i_m_axis_rx_tdata[13: 12];
                    v.req_len = i_m_axis_rx_tdata[9: 0];
                    v.req_rid = i_m_axis_rx_tdata[63: 48];
                    v.req_tag = i_m_axis_rx_tdata[47: 40];
                    v.req_be = i_m_axis_rx_tdata[39: 32];
                    v.state = PIO_RX_MEM_RD32_DW1DW2;
                end else begin
                    v.state = PIO_RX_RST_STATE;
                end
            end

            PIO_RX_MEM_WR32_FMT_TYPE: begin
                if (i_m_axis_rx_tdata[9: 0] == 10'd1) begin
                    v.wr_be = i_m_axis_rx_tdata[39: 32];
                    v.state = PIO_RX_MEM_WR32_DW1DW2;
                end else begin
                    v.state = PIO_RX_RST_STATE;
                end
            end

            PIO_RX_MEM_RD64_FMT_TYPE: begin
                if (i_m_axis_rx_tdata[9: 0] == 10'd1) begin
                    v.req_tc = i_m_axis_rx_tdata[22: 20];
                    v.req_td = i_m_axis_rx_tdata[15];
                    v.req_ep = i_m_axis_rx_tdata[14];
                    v.req_attr = i_m_axis_rx_tdata[13: 12];
                    v.req_len = i_m_axis_rx_tdata[9: 0];
                    v.req_rid = i_m_axis_rx_tdata[63: 48];
                    v.req_tag = i_m_axis_rx_tdata[47: 40];
                    v.req_be = i_m_axis_rx_tdata[39: 32];
                    v.state = PIO_RX_MEM_RD64_DW1DW2;
                end else begin
                    v.state = PIO_RX_RST_STATE;
                end
            end

            PIO_RX_MEM_WR64_FMT_TYPE: begin
                if (i_m_axis_rx_tdata[9: 0] == 10'd1) begin
                    v.wr_be = i_m_axis_rx_tdata[39: 32];
                    v.state = PIO_RX_MEM_WR64_DW1DW2;
                end else begin
                    v.state = PIO_RX_RST_STATE;
                end
            end

            PIO_RX_IO_RD32_FMT_TYPE: begin
                if (i_m_axis_rx_tdata[9: 0] == 10'd1) begin
                    v.req_tc = i_m_axis_rx_tdata[22: 20];
                    v.req_td = i_m_axis_rx_tdata[15];
                    v.req_ep = i_m_axis_rx_tdata[14];
                    v.req_attr = i_m_axis_rx_tdata[13: 12];
                    v.req_len = i_m_axis_rx_tdata[9: 0];
                    v.req_rid = i_m_axis_rx_tdata[63: 48];
                    v.req_tag = i_m_axis_rx_tdata[47: 40];
                    v.req_be = i_m_axis_rx_tdata[39: 32];
                    v.state = PIO_RX_MEM_RD32_DW1DW2;
                end else begin
                    v.state = PIO_RX_RST_STATE;
                end
            end

            PIO_RX_IO_WR32_FMT_TYPE: begin
                if (i_m_axis_rx_tdata[9: 0] == 10'd1) begin
                    v.req_tc = i_m_axis_rx_tdata[22: 20];
                    v.req_td = i_m_axis_rx_tdata[15];
                    v.req_ep = i_m_axis_rx_tdata[14];
                    v.req_attr = i_m_axis_rx_tdata[13: 12];
                    v.req_len = i_m_axis_rx_tdata[9: 0];
                    v.req_rid = i_m_axis_rx_tdata[63: 48];
                    v.req_tag = i_m_axis_rx_tdata[47: 40];
                    v.req_be = i_m_axis_rx_tdata[39: 32];
                    v.wr_be = i_m_axis_rx_tdata[39: 32];
                    v.state = PIO_RX_IO_WR_DW1DW2;
                end else begin
                    v.state = PIO_RX_RST_STATE;
                end
            end

            default: begin
                v.state = PIO_RX_RST_STATE;
            end
            endcase
        end else begin
            v.state = PIO_RX_RST_STATE;
        end
    end

    PIO_RX_MEM_RD32_DW1DW2: begin
        if (i_m_axis_rx_tvalid == 1'b1) begin
            v.m_axis_rx_tready = 1'b0;
            v.req_valid = 1'b1;
            v.req_addr = {vb_region_select[1: 0], i_m_axis_rx_tdata[10: 2], 2'd0};
            v.tlp_resp = TLP_POSTED;
            v.state = PIO_RX_WAIT_DMA_RESP;
        end else begin
            v.state = PIO_RX_MEM_RD32_DW1DW2;
        end
    end

    PIO_RX_MEM_WR32_DW1DW2: begin
        if (i_m_axis_rx_tvalid == 1'b1) begin
            v.m_axis_rx_tready = 1'b0;
            v.req_valid = 1'b1;
            v.wr_en = 1'b1;
            v.wr_addr = {vb_region_select[1: 0], i_m_axis_rx_tdata[10: 2]};
            v.req_addr = {vb_region_select[1: 0], i_m_axis_rx_tdata[10: 2], 2'd0};
            v.wr_data = {i_m_axis_rx_tdata[63: 32], i_m_axis_rx_tdata[63: 32]};
            if (i_m_axis_rx_tdata[2] == 1'b1) begin
                v.wr_be = {r.wr_be[3: 0], r.wr_be[7: 4]};
            end
            v.tlp_resp = TLP_NON_POSTED;
            v.state = PIO_RX_WAIT_DMA_RESP;
        end else begin
            v.state = PIO_RX_MEM_WR32_DW1DW2;
        end
    end

    PIO_RX_MEM_RD64_DW1DW2: begin
        if (i_m_axis_rx_tvalid == 1'b1) begin
            v.m_axis_rx_tready = 1'b0;
            v.req_valid = 1'b1;
            v.req_addr = {vb_region_select[1: 0], i_m_axis_rx_tdata[42: 34], 2'd0};
            v.tlp_resp = TLP_POSTED;
            v.state = PIO_RX_WAIT_DMA_RESP;
        end else begin
            v.state = PIO_RX_MEM_RD64_DW1DW2;
        end
    end

    PIO_RX_MEM_WR64_DW1DW2: begin
        if (i_m_axis_rx_tvalid == 1'b1) begin
            v.wr_addr = {vb_region_select[1: 0], i_m_axis_rx_tdata[42: 34]};
            v.req_addr = {vb_region_select[1: 0], i_m_axis_rx_tdata[42: 34], 2'd0};
            if (i_m_axis_rx_tdata[34] == 1'b1) begin
                v.wr_be = {r.wr_be[3: 0], r.wr_be[7: 4]};
            end
            v.state = PIO_RX_MEM_WR64_DW3;
        end else begin
            v.state = PIO_RX_MEM_WR64_DW1DW2;
        end
    end

    PIO_RX_MEM_WR64_DW3: begin
        if (i_m_axis_rx_tvalid == 1'b1) begin
            v.m_axis_rx_tready = 1'b0;
            v.req_valid = 1'b1;
            v.wr_en = 1'b1;
            v.wr_data = {i_m_axis_rx_tdata[31: 0], i_m_axis_rx_tdata[31: 0]};
            v.tlp_resp = TLP_NON_POSTED;
            v.state = PIO_RX_WAIT_DMA_RESP;
        end else begin
            v.state = PIO_RX_MEM_WR64_DW3;
        end
    end

    PIO_RX_IO_WR_DW1DW2: begin
        if (i_m_axis_rx_tvalid == 1'b1) begin
            v.m_axis_rx_tready = 1'b0;
            v.req_valid = 1'b1;
            v.wr_en = 1'b1;
            v.wr_addr = {vb_region_select[1: 0], i_m_axis_rx_tdata[10: 2]};
            v.req_addr = {vb_region_select[1: 0], i_m_axis_rx_tdata[10: 2], 2'd0};
            v.wr_data = {i_m_axis_rx_tdata[63: 32], i_m_axis_rx_tdata[63: 32]};
            if (i_m_axis_rx_tdata[2] == 1'b1) begin
                v.wr_be = {r.wr_be[3: 0], r.wr_be[7: 4]};
            end
            v.tlp_resp = TLP_COMPLETION;
            v.state = PIO_RX_WAIT_DMA_RESP;
        end else begin
            v.state = PIO_RX_IO_WR_DW1DW2;
        end
    end

    PIO_RX_WAIT_DMA_RESP: begin
        if (i_req_mem_ready == 1'b1) begin
            v.req_valid = 1'b0;
        end
        if (i_resp_mem_valid == 1'b1) begin
            if ((|r.tlp_resp) == 1'b1) begin
                v.tlp_resp = 2'd0;
                v.state = PIO_RX_WAIT_TX_COMPLETION;
            end else begin
                v.m_axis_rx_tready = 1'b1;
                v.state = PIO_RX_RST_STATE;
            end
        end
    end

    PIO_RX_WAIT_TX_COMPLETION: begin
        v.wr_en = 1'b0;
        v.req_len = 10'd0;
        if (i_compl_done == 1'b1) begin
            v.m_axis_rx_tready = 1'b1;
            v.state = PIO_RX_RST_STATE;
        end
    end

    default: begin
        v.state = PIO_RX_RST_STATE;
    end
    endcase

    rin = v;
end: comb_proc


assign o_m_axis_rx_tready = r.m_axis_rx_tready;
assign o_req_compl = r.tlp_resp[0];
assign o_req_compl_wd = r.tlp_resp[1];
assign o_req_tc = r.req_tc;
assign o_req_td = r.req_td;
assign o_req_ep = r.req_ep;
assign o_req_attr = r.req_attr;
assign o_req_len = r.req_len;
assign o_req_rid = r.req_rid;
assign o_req_tag = r.req_tag;
assign o_req_be = r.req_be;
assign o_req_addr = r.req_addr;

assign o_req_mem_valid = r.req_valid;
assign o_req_mem_64 = 1'b0;
assign o_req_mem_write = r.wr_en;
assign o_req_mem_bytes = {r.req_len, 2'd0};
assign o_req_mem_addr = r.req_addr;
assign o_req_mem_strob = r.wr_be;
assign o_req_mem_data = r.wr_data;
assign o_req_mem_last = 1'b1;

always_ff @(posedge i_clk, negedge i_nrst) begin
    if (i_nrst == 1'b0) begin
        r <= pcie_io_rx_engine_r_reset;
    end else begin
        r <= rin;
    end
end

endmodule: pcie_io_rx_engine
