// 
//  Copyright 2022 Sergey Khabarov, sergeykhbr@gmail.com
// 
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
// 

`timescale 1ns/10ps

module pcie_dma #(
    parameter bit async_reset = 1'b0
)
(
    input logic i_nrst,                                     // System Reset: active LOW
    input logic i_clk,                                      // System bus clock
    input logic i_pcie_phy_clk,                             // PCIE clock generated by end-point
    // PCIE EP - DMA engine interface
    input logic [15:0] i_pcie_completer_id,                 // Bus, Device, Function
    output logic [3:0] o_dma_state,                         // State machine debug output, connected to APB controller
    input types_dma_pkg::pcie_dma64_in_type i_pcie_dmai,    // PCIE-EP to system DMA requests
    output types_dma_pkg::pcie_dma64_out_type o_pcie_dmao,  // System DMA responds to PCIE EP
    // DMA engine interface - System on Chip interface
    output types_pnp_pkg::dev_config_type o_xmst_cfg,       // PCIE DMA master interface descriptor
    input types_amba_pkg::axi4_master_in_type i_xmsti,
    output types_amba_pkg::axi4_master_out_type o_xmsto
);

import types_dma_pkg::*;
import types_pnp_pkg::*;
import types_amba_pkg::*;
import pcie_cfg_pkg::*;
import pcie_dma_pkg::*;

logic [REQ_FIFO_WIDTH-1:0] wb_reqfifo_payload_i;
logic [REQ_FIFO_WIDTH-1:0] wb_reqfifo_payload_o;
logic w_reqfifo_full;
logic w_reqfifo_empty;
logic w_reqfifo_rd;
logic [RESP_FIFO_WIDTH-1:0] wb_respfifo_payload_i;
logic [RESP_FIFO_WIDTH-1:0] wb_respfifo_payload_o;
logic w_respfifo_full;
logic w_respfifo_empty;
logic w_respfifo_wr;
pcie_dma_registers r, rin;

// PCIE EP (200 MHz) -> DMA (40 MHz)
cdc_afifo #(
    .abits(CFG_PCIE_DMAFIFO_DEPTH),
    .dbits(REQ_FIFO_WIDTH)
) reqfifo (
    .i_nrst(i_nrst),
    .i_wclk(i_pcie_phy_clk),
    .i_wr(i_pcie_dmai.valid),
    .i_wdata(wb_reqfifo_payload_i),
    .o_wfull(w_reqfifo_full),
    .i_rclk(i_clk),
    .i_rd(w_reqfifo_rd),
    .o_rdata(wb_reqfifo_payload_o),
    .o_rempty(w_reqfifo_empty)
);
// DMA (40 MHz) -> PCIE EP (200 MHz)
cdc_afifo #(
    .abits(CFG_PCIE_DMAFIFO_DEPTH),
    .dbits(RESP_FIFO_WIDTH)
) respfifo (
    .i_nrst(i_nrst),
    .i_wclk(i_clk),
    .i_wr(w_respfifo_wr),
    .i_wdata(wb_respfifo_payload_i),
    .o_wfull(w_respfifo_full),
    .i_rclk(i_pcie_phy_clk),
    .i_rd(i_pcie_dmai.ready),
    .o_rdata(wb_respfifo_payload_o),
    .o_rempty(w_respfifo_empty)
);

always_comb
begin: comb_proc
    pcie_dma_registers v;
    dev_config_type vb_xmst_cfg;
    axi4_master_out_type vb_xmsto;
    logic [XSIZE_TOTAL-1:0] vb_xbytes;                      // result of function call XSize2XBytes(xsize)
    logic v_req_ready;
    logic [63:0] vb_req_addr;
    logic [1:0] vb_req_addr1_0;                             // address[1:0] restored from strob field be[3:0]
    logic [63:0] vb_req_data;
    logic [7:0] vb_req_strob;
    logic v_req_last;
    logic v_single_tlp;                                     // single 32-bit dma transaction, trnasmit as 4DW with TLP header
    logic v_resp_valid;
    logic [63:0] vb_resp_data;
    logic [7:0] vb_resp_strob;
    logic v_resp_last;

    vb_xmst_cfg = dev_config_none;
    vb_xmsto = axi4_master_out_none;
    vb_xbytes = 8'd0;
    v_req_ready = 1'b0;
    vb_req_addr = 64'd0;
    vb_req_addr1_0 = 2'd0;
    vb_req_data = 64'd0;
    vb_req_strob = 8'd0;
    v_req_last = 1'b0;
    v_single_tlp = 1'b0;
    v_resp_valid = 1'b0;
    vb_resp_data = 64'd0;
    vb_resp_strob = 8'd0;
    v_resp_last = 1'b0;

    v = r;

    v_req_ready = 1'b0;
    vb_req_addr = 64'd0;
    v_resp_valid = 1'b0;
    vb_resp_data = 64'd0;
    vb_resp_strob = 8'd0;
    v_resp_last = 1'b0;
    v_single_tlp = 1'b0;
    vb_xmsto = axi4_master_out_none;

    if (r.dw0[9: 0] == 10'd1) begin
        // DW0[9:0] = Length number of DW (4-bytes) for 32/64 bars
        v_single_tlp = 1'b1;
    end
    vb_xmst_cfg.descrsize = PNP_CFG_DEV_DESCR_BYTES;
    vb_xmst_cfg.descrtype = PNP_CFG_TYPE_MASTER;
    vb_xmst_cfg.vid = VENDOR_OPTIMITECH;
    vb_xmst_cfg.did = OPTIMITECH_PCIE_DMA;
    vb_xbytes = XSizeToBytes(r.xsize);

    // Request address bits [1:0] are not transmitted, should be restored from BE[3:0]:
    // be[3:0] => addr[1:0]
    // 0000    => 00
    // xxx1    => 00
    // xx10    => 01
    // x100    => 10
    // 1000    => 11
    if (r.dw1[0] == 1'b1) begin
        vb_req_addr1_0 = 2'd0;
    end else if (r.dw1[1] == 1'b1) begin
        vb_req_addr1_0 = 2'd1;
    end else if (r.dw1[2] == 1'b1) begin
        vb_req_addr1_0 = 2'd2;
    end else if (r.dw1[3] == 1'b1) begin
        vb_req_addr1_0 = 2'd3;
    end else begin
        vb_req_addr1_0 = 2'd0;
    end

    // Request FIFO inputs/outputs:
    wb_reqfifo_payload_i = {i_pcie_dmai.last,
            i_pcie_dmai.strob,
            i_pcie_dmai.data};

    v_req_last = wb_reqfifo_payload_o[72];
    vb_req_strob = wb_reqfifo_payload_o[71: 64];
    vb_req_data = wb_reqfifo_payload_o[63: 0];

    // Temporary register
    case (r.state)
    STATE_RST: begin
        v_req_ready = 1'b1;
        v.resp_status = TLP_STATUS_SUCCESS;
        v.req_rd_locked = 1'b0;
        v.resp_cpl = 7'd0;
        v.resp_with_payload = 1'b0;
        if (w_reqfifo_empty == 1'b0) begin
            v.dw0 = vb_req_data[31: 0];
            v.dw1 = vb_req_data[63: 32];
            v.state = STATE_DW3DW4;
        end
    end

    STATE_DW3DW4: begin
        // 64-bits BAR could use 3DW header because if addr[63:32] is zero
        // TLP behaviour is undefined (Xilinx example ignores it):
        //   dw2 = addr[63:32]
        //   dw3 = {addr[31:2], 00}
        v_req_ready = 1'b1;
        v.xlen = (r.dw0[7: 0] - 1);                         // warning: Actual size of Length is 10 bits. 0 is 1024 DWs (4096 Bytes)
        v.dw2 = vb_req_data[31: 0];
        v.dw3 = 32'd0;
        if (w_reqfifo_empty == 1'b0) begin
            // fmt[0] = 1 when 4DW header is used
            if (r.dw0[29] == 1'b1) begin
                v.dw3 = vb_req_data[63: 32];
            end
            if (r.dw0[30] == 1'b0) begin
                // fmt[1]=0: read operation
                v.state = STATE_AR;
                case (r.dw0[28: 24])                        // DW0[28:24] = Type[4:0]
                5'h01: begin
                    // Read Locked request (in case of error becomes PCIE_CPL_LOCKED_READ_NODATA:
                    v.resp_cpl = PCIE_CPL_LOCKED_READ;
                    v.req_rd_locked = 1'b1;
                end
                5'h02: begin
                    // I/O Read request:
                    v.resp_cpl = PCIE_CPL_DATA;
                end
                5'h05: begin
                    // Configuration Read request Root Port (type 1):
                    v.resp_cpl = PCIE_CPL_DATA;
                end
                default: begin
                    // Read request.
                    v.resp_cpl = PCIE_CPL_DATA;
                end
                endcase

                v.byte_cnt = {r.dw0[7: 0], 2'd0};
                if (r.dw0[29] == 1'b0) begin
                    // fmt[0]=0: 3DW header (32-bits address):
                    v.xsize = 3'd2;
                    vb_req_addr[31: 0] = {vb_req_data[31: 2], vb_req_addr1_0};
                end else begin
                    // fmt[0]=1: 4DW header (64-bits address):
                    v.xsize = 3'd3;
                    vb_req_addr = {vb_req_data[31: 0], vb_req_data[63: 34], vb_req_addr1_0};
                end
            end else begin
                // fmt[1] = 1: write operation
                v.state = STATE_AW;
                v.xwstrb = r.dw1[7: 0];
                case (r.dw0[28: 24])                        // DW0[28:24] = Type[4:0]
                5'h02: begin
                    // I/O Write request:
                    v.resp_cpl = PCIE_CPL_NODATA;
                end
                5'h05: begin
                    // Configuration Write request Root Port (type 1):
                    v.resp_cpl = PCIE_CPL_NODATA;
                end
                default: begin
                    // Write request. No completion.
                end
                endcase

                v.byte_cnt = {r.dw0[7: 0], 2'd0};
                if (r.dw0[29] == 1'b0) begin
                    // fmt[0]=0: 3DW header (32-bits address):
                    v.xsize = 3'd2;
                    vb_req_addr[31: 0] = {vb_req_data[31: 2], vb_req_addr1_0};
                    v.xwdata = {vb_req_data[63: 32], vb_req_data[63: 32]};
                    v.xwena = v_req_last;                   // AXI Light: burst transactions are no supported
                end else begin
                    // fmt[0]=1: 4DW header (64-bits address):
                    v.xsize = 3'd3;
                    vb_req_addr = {vb_req_data[31: 0], vb_req_data[63: 34], vb_req_addr1_0};
                end
            end
        end
        v.xaddr = vb_req_addr[(CFG_SYSBUS_ADDR_BITS - 1): 0];
    end
    STATE_AR: begin
        vb_xmsto.ar_valid = 1'b1;
        vb_xmsto.ar_bits.addr = r.xaddr[(CFG_SYSBUS_ADDR_BITS - 1): 0];
        // sram base address: 64'h0000000008000000
        vb_xmsto.ar_bits.addr = {36'h000008001, vb_xmsto.ar_bits.addr[11: 0]};
        vb_xmsto.ar_bits.len = r.xlen;
        vb_xmsto.ar_bits.size = r.xsize;
        vb_xmsto.ar_bits.lock = r.req_rd_locked;
        v.resp_with_payload = 1'b1;
        if (i_xmsti.ar_ready == 1'b1) begin
            if (v_single_tlp == 1'b1) begin
                // 3DW header + DW 32-bits payload
                v.state = STATE_R_SINGLE32;
            end else begin
                // 3DW header only
                v.state = STATE_RESP_DW0DW1;
            end
        end
    end
    STATE_R_SINGLE32: begin
        // 32-bit single transactions (no bulk). MEM32 and IO only:
        vb_xmsto.r_ready = 1'b1;
        v.xerr = i_xmsti.r_resp;
        if (r.xaddr[2] == 1'b0) begin
            v.xrdata = {i_xmsti.r_data[31: 0], i_xmsti.r_data[31: 0]};
        end else begin
            v.xrdata = {i_xmsti.r_data[63: 32], i_xmsti.r_data[63: 32]};
        end
        if (i_xmsti.r_valid == 1'b1) begin
            v.state = STATE_RESP_DW0DW1;
        end
    end
    STATE_R: begin
        vb_xmsto.r_ready = (~w_reqfifo_full);
        v_resp_valid = i_xmsti.r_valid;
        vb_resp_strob = 8'hFF;
        v_resp_last = (~(|r.xlen));
        v.xerr = i_xmsti.r_resp;
        if (r.xsize == 3'd2) begin
            // 32-bit transactions:
            if (r.xaddr[2] == 1'b0) begin
                vb_resp_data = {i_xmsti.r_data[31: 0], i_xmsti.r_data[31: 0]};
            end else begin
                vb_resp_data = {i_xmsti.r_data[63: 32], i_xmsti.r_data[63: 32]};
            end
        end else begin
            // 64-bit transactions:
            vb_resp_data = i_xmsti.r_data;
        end

        if ((i_xmsti.r_valid == 1'b1) && (w_respfifo_full == 1'b0)) begin
            // Burst support: 
            if (i_xmsti.r_resp != AXI_RESP_OKAY) begin
                v.resp_status = TLP_STATUS_ABORTED;
                if (r.req_rd_locked == 1'b1) begin
                    // Error on Locked Read transaction:
                    v.resp_cpl = PCIE_CPL_LOCKED_READ_NODATA;
                end
                v.state = STATE_RESP_DW0DW1;
            end else if ((|r.xlen) == 1'b1) begin
                v.xlen = (r.xlen - 1);
                v.xaddr = (r.xaddr + vb_xbytes);
                v.byte_cnt = (r.byte_cnt - vb_xbytes);
            end else begin
                v.state = STATE_RST;
            end
        end
    end
    STATE_AW: begin
        vb_xmsto.aw_valid = 1'b1;
        vb_xmsto.aw_bits.addr = r.xaddr[(CFG_SYSBUS_ADDR_BITS - 1): 0];
        // sram base address: 64'h0000000008000000
        vb_xmsto.aw_bits.addr = {36'h000008001, vb_xmsto.aw_bits.addr[11: 0]};
        vb_xmsto.aw_bits.len = r.xlen;
        vb_xmsto.aw_bits.size = r.xsize;
        vb_xmsto.w_valid = r.xwena;
        vb_xmsto.w_last = r.xwena;
        vb_xmsto.w_strb = r.xwstrb;
        vb_xmsto.w_data = {r.xwdata[31: 0], r.xwdata[31: 0]};
        if (i_xmsti.aw_ready == 1'b1) begin
            if ((r.xwena == 1'b1) && (i_xmsti.w_ready == 1'b1)) begin
                // AXI light: no burst transactions:
                v.state = STATE_B;
                v.xwena = 1'b0;
            end else begin
                v.state = STATE_W;
            end
        end
    end
    STATE_W: begin
        if (r.xwena == 1'b1) begin
            v.xwena = 1'b0;
            vb_xmsto.w_valid = 1'b1;
            vb_xmsto.w_strb = r.xwstrb;
            vb_xmsto.w_data = r.xwdata;
            vb_xmsto.w_last = 1'b1;
            if (i_xmsti.w_ready == 1'b1) begin
                v.state = STATE_B;
            end
        end else begin
            v_req_ready = i_xmsti.w_ready;
            vb_xmsto.w_valid = (~w_reqfifo_empty);
            vb_xmsto.w_strb = vb_req_strob;
            vb_xmsto.w_data = vb_req_data;
            vb_xmsto.w_last = (~(|r.xlen));
            if ((w_reqfifo_empty == 1'b0) && (i_xmsti.w_ready == 1'b1)) begin
                if (v_req_last == 1'b1) begin
                    v.state = STATE_B;
                end
            end
        end
    end
    STATE_B: begin
        vb_xmsto.b_ready = 1'b1;
        if (i_xmsti.b_valid == 1'b1) begin
            v.xerr = i_xmsti.b_resp;
            if (i_xmsti.b_resp != AXI_RESP_OKAY) begin
                v.resp_status = TLP_STATUS_ABORTED;
            end
            if ((|r.resp_cpl) == 1'b0) begin
                // Posted write TLP without response
                v.state = STATE_RST;
            end else begin
                // Non-posted write TLP with response
                v.state = STATE_RESP_DW0DW1;
            end
        end
    end

    STATE_RESP_DW0DW1: begin
        v_resp_valid = 1'b1;
        vb_resp_strob = 8'hFF;
        vb_resp_data[9: 0] = r.dw0[9: 0];                   // DW0[9:0] Length
        vb_resp_data[11: 10] = 2'd0;                        // DW0[11:10] Reserved
        vb_resp_data[13: 12] = r.dw0[13: 12];               // DW0[13:12] Attr
        vb_resp_data[14] = r.dw0[14];                       // DW0[14] EP
        vb_resp_data[15] = r.dw0[15];                       // DW0[15] TD
        vb_resp_data[19: 16] = 4'd0;                        // DW0[19:16] Reserved
        vb_resp_data[22: 20] = r.dw0[22: 20];               // DW0[22:20] TC
        vb_resp_data[23] = 1'b0;                            // DW0[23] Reserved
        vb_resp_data[30: 24] = r.resp_cpl;                  // DW0[30:24] {Fmt,Type} Completion
        vb_resp_data[31] = 1'b0;                            // DW0[31] Reserved
        vb_resp_data[43: 32] = r.byte_cnt;                  // DW1[11:0] Byte Count
        vb_resp_data[44] = 1'b0;                            // DW1[12] BCM
        vb_resp_data[47: 45] = r.resp_status;               // DW1[15:13] Status
        vb_resp_data[63: 48] = i_pcie_completer_id;         // DW1[31:16] Completer ID
        if (w_respfifo_full == 1'b0) begin
            v.state = STATE_RESP_DW2DW3;
        end
    end

    STATE_RESP_DW2DW3: begin
        v_resp_valid = 1'b1;
        vb_resp_strob = 8'h0F;
        vb_resp_data[6: 0] = r.xaddr[6: 0];                 // DW2[6:0] Low Address
        vb_resp_data[7] = 1'b0;                             // DW2[7] Reserved
        vb_resp_data[15: 8] = r.dw1[15: 8];                 // DW2[15:8] Tag
        vb_resp_data[31: 16] = r.dw1[31: 16];               // DW2[31:16] Requester ID
        vb_resp_data[63: 32] = r.xrdata[31: 0];             // DW3[31:0] payload (ignored by strob 0F)
        if (w_respfifo_full == 1'b0) begin
            if (r.resp_status != TLP_STATUS_SUCCESS) begin
                v_resp_last = 1'b1;
                v.state = STATE_RST;
            end else if ((v_single_tlp == 1'b1) && (r.resp_with_payload == 1'b1)) begin
                // DW4 response with the single DW payload
                vb_resp_strob = 8'hFF;
                v_resp_last = 1'b1;
                v.state = STATE_RST;
            end else if (r.resp_with_payload == 1'b1) begin
                // DW3 response only if: payload not a single tlp32
                v.state = STATE_R;
            end else begin
                // DW3 without payload
                v_resp_last = 1'b1;
                v.state = STATE_RST;
            end
        end
    end

    default: begin
        v.state = STATE_RST;
    end
    endcase

    if (~async_reset && i_nrst == 1'b0) begin
        v = pcie_dma_r_reset;
    end

    // Response FIFO inputs/outputs:
    wb_respfifo_payload_i = {v_resp_last,
            vb_resp_strob,
            vb_resp_data};
    o_pcie_dmao.last = wb_respfifo_payload_o[72];
    o_pcie_dmao.strob = wb_respfifo_payload_o[71: 64];
    o_pcie_dmao.data = wb_respfifo_payload_o[63: 0];
    o_pcie_dmao.ready = (~w_reqfifo_full);
    o_pcie_dmao.valid = (~w_respfifo_empty);
    w_respfifo_wr = v_resp_valid;
    w_reqfifo_rd = v_req_ready;
    o_xmst_cfg = vb_xmst_cfg;
    o_xmsto = vb_xmsto;

    rin = v;
end: comb_proc


generate
    if (async_reset) begin: async_rst_gen

        always_ff @(posedge i_clk, negedge i_nrst) begin: rg_proc
            if (i_nrst == 1'b0) begin
                r <= pcie_dma_r_reset;
            end else begin
                r <= rin;
            end
        end: rg_proc

    end: async_rst_gen
    else begin: no_rst_gen

        always_ff @(posedge i_clk) begin: rg_proc
            r <= rin;
        end: rg_proc

    end: no_rst_gen
endgenerate

endmodule: pcie_dma
