// 
//  Copyright 2022 Sergey Khabarov, sergeykhbr@gmail.com
// 
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
// 

`timescale 1ns/10ps

module pcie_dma(
    input logic i_nrst,                                     // System Reset: active LOW
    input logic i_clk,                                      // System bus clock
    input logic i_pcie_phy_clk,                             // PCIE clock generated by end-point
    // PCIE EP - DMA engine interface
    input logic [15:0] i_pcie_completer_id,                 // Bus, Device, Function
    output logic [3:0] o_dma_state,                         // State machine debug output, connected to APB controller
    input types_dma_pkg::pcie_dma64_in_type i_pcie_dmai,    // PCIE-EP to system DMA requests
    output types_dma_pkg::pcie_dma64_out_type o_pcie_dmao,  // System DMA responds to PCIE EP
    // DMA engine interface - System on Chip interface
    output types_pnp_pkg::dev_config_type o_xmst_cfg,       // PCIE DMA master interface descriptor
    input types_amba_pkg::axi4_master_in_type i_xmsti,
    output types_amba_pkg::axi4_master_out_type o_xmsto,
    // Debug signals:
    output logic o_dbg_mem_valid,
    output logic o_dbg_mem_wren,
    output logic [7:0] o_dbg_mem_wstrb,
    output logic [12:0] o_dbg_mem_addr,
    output logic [31:0] o_dbg_mem_data
);

import types_dma_pkg::*;
import types_pnp_pkg::*;
import types_amba_pkg::*;
import pcie_cfg_pkg::*;
import pcie_dma_pkg::*;

logic w_pcie_dmai_valid;
logic w_pcie_dmai_ready;
logic [REQ_FIFO_WIDTH-1:0] wb_reqfifo_payload_i;
logic [REQ_FIFO_WIDTH-1:0] wb_reqfifo_payload_o;
logic w_reqfifo_wready;
logic w_reqfifo_rvalid;
logic w_reqfifo_rd;
logic [RESP_FIFO_WIDTH-1:0] wb_respfifo_payload_i;
logic [RESP_FIFO_WIDTH-1:0] wb_respfifo_payload_o;
logic w_respfifo_wready;
logic w_respfifo_rvalid;
logic w_respfifo_wr;
logic [8:0] wb_m_axis_rx_tuser;
logic w_m_axis_rx_tlast;
logic [KEEP_WIDTH-1:0] wb_m_axis_rx_tkeep;
logic [C_DATA_WIDTH-1:0] wb_m_axis_rx_tdata;
logic w_s_axis_tx_tlast;
logic [KEEP_WIDTH-1:0] wb_s_axis_tx_tkeep;
logic [C_DATA_WIDTH-1:0] wb_s_axis_tx_tdata;
logic w_tx_src_dsc;
logic w_req_compl;
logic w_compl_done;

// PCIE EP (200 MHz) -> DMA (40 MHz)
cdc_afifo #(
    .abits(CFG_PCIE_DMAFIFO_DEPTH),
    .dbits(REQ_FIFO_WIDTH)
) reqfifo (
    .i_nrst(i_nrst),
    .i_wclk(i_pcie_phy_clk),
    .i_wr(w_pcie_dmai_valid),
    .i_wdata(wb_reqfifo_payload_i),
    .o_wready(w_reqfifo_wready),
    .i_rclk(i_clk),
    .i_rd(w_reqfifo_rd),
    .o_rdata(wb_reqfifo_payload_o),
    .o_rvalid(w_reqfifo_rvalid)
);
// DMA (40 MHz) -> PCIE EP (200 MHz)
cdc_afifo #(
    .abits(CFG_PCIE_DMAFIFO_DEPTH),
    .dbits(RESP_FIFO_WIDTH)
) respfifo (
    .i_nrst(i_nrst),
    .i_wclk(i_clk),
    .i_wr(w_respfifo_wr),
    .i_wdata(wb_respfifo_payload_i),
    .o_wready(w_respfifo_wready),
    .i_rclk(i_pcie_phy_clk),
    .i_rd(w_pcie_dmai_ready),
    .o_rdata(wb_respfifo_payload_o),
    .o_rvalid(w_respfifo_rvalid)
);

pcie_io_ep #(
    .C_DATA_WIDTH(C_DATA_WIDTH),
    .KEEP_WIDTH(KEEP_WIDTH)
) PIO_EP_inst (
    .i_nrst(i_nrst),
    .i_clk(i_clk),
    .i_s_axis_tx_tready(w_respfifo_wready),
    .o_s_axis_tx_tdata(wb_s_axis_tx_tdata),
    .o_s_axis_tx_tkeep(wb_s_axis_tx_tkeep),
    .o_s_axis_tx_tlast(w_s_axis_tx_tlast),
    .o_s_axis_tx_tvalid(w_respfifo_wr),
    .o_tx_src_dsc(w_tx_src_dsc),
    .i_m_axis_rx_tdata(wb_m_axis_rx_tdata),
    .i_m_axis_rx_tkeep(wb_m_axis_rx_tkeep),
    .i_m_axis_rx_tlast(w_m_axis_rx_tlast),
    .i_m_axis_rx_tvalid(w_reqfifo_rvalid),
    .o_m_axis_rx_tready(w_reqfifo_rd),
    .i_m_axis_rx_tuser(wb_m_axis_rx_tuser),
    .o_req_compl(w_req_compl),
    .o_compl_done(w_compl_done),
    .i_cfg_completer_id(i_pcie_completer_id),
    .o_mem_valid(o_dbg_mem_valid),
    .o_mem_wren(o_dbg_mem_wren),
    .o_mem_wstrb(o_dbg_mem_wstrb),
    .o_mem_addr(o_dbg_mem_addr),
    .o_mem_data(o_dbg_mem_data)
);

always_comb
begin: comb_proc
    dev_config_type vb_xmst_cfg;
    axi4_master_out_type vb_xmsto;
    pcie_dma64_out_type vb_pcie_dmao;
    logic [8:0] vb_m_axis_rx_tuser;
    logic v_m_axis_rx_tlast;
    logic [KEEP_WIDTH-1:0] vb_m_axis_rx_tkeep;
    logic [C_DATA_WIDTH-1:0] vb_m_axis_rx_tdata;

    vb_m_axis_rx_tuser = 9'd0;
    v_m_axis_rx_tlast = 1'b0;
    vb_m_axis_rx_tkeep = 8'd0;
    vb_m_axis_rx_tdata = 64'd0;

    vb_xmst_cfg.descrsize = PNP_CFG_DEV_DESCR_BYTES;
    vb_xmst_cfg.descrtype = PNP_CFG_TYPE_MASTER;
    vb_xmst_cfg.vid = VENDOR_OPTIMITECH;
    vb_xmst_cfg.did = OPTIMITECH_PCIE_DMA;
    o_xmst_cfg = vb_xmst_cfg;
    o_xmsto = axi4_master_out_none;

    o_dma_state = '0;

    // PCIE PHY clock to system clock AFIFO:

    // SystemC limitation, cannot assign directly to signal:
    vb_m_axis_rx_tuser = wb_reqfifo_payload_o[81: 73];
    v_m_axis_rx_tlast = wb_reqfifo_payload_o[72];
    vb_m_axis_rx_tkeep = wb_reqfifo_payload_o[71: 64];
    vb_m_axis_rx_tdata = wb_reqfifo_payload_o[63: 0];
    wb_m_axis_rx_tuser = vb_m_axis_rx_tuser;
    w_m_axis_rx_tlast = v_m_axis_rx_tlast;
    wb_m_axis_rx_tkeep = vb_m_axis_rx_tkeep;
    wb_m_axis_rx_tdata = vb_m_axis_rx_tdata;

    vb_pcie_dmao.valid = w_respfifo_rvalid;
    vb_pcie_dmao.ready = w_reqfifo_wready;
    vb_pcie_dmao.last = wb_respfifo_payload_o[72];
    vb_pcie_dmao.strob = wb_respfifo_payload_o[71: 64];
    vb_pcie_dmao.data = wb_respfifo_payload_o[63: 0];
    o_pcie_dmao = vb_pcie_dmao;
end: comb_proc


assign w_pcie_dmai_valid = i_pcie_dmai.valid;
assign w_pcie_dmai_ready = i_pcie_dmai.ready;
assign wb_reqfifo_payload_i = {i_pcie_dmai.bar_hit,
        i_pcie_dmai.ecrc_err,
        i_pcie_dmai.err_fwd,
        i_pcie_dmai.last,
        i_pcie_dmai.strob,
        i_pcie_dmai.data};

// System Clock to PCIE PHY clock AFIFO:
assign wb_respfifo_payload_i = {w_s_axis_tx_tlast,
        wb_s_axis_tx_tkeep,
        wb_s_axis_tx_tdata};

endmodule: pcie_dma
