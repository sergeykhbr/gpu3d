// 
//  Copyright 2022 Sergey Khabarov, sergeykhbr@gmail.com
// 
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
// 

`timescale 1ns/10ps

module pcie_dma(
    input logic i_sys_nrst,                                 // System Reset: active LOW
    input logic i_sys_clk,                                  // System bus clock
    input logic i_pcie_usr_rst,                             // PCIE user rest: active HIGH
    input logic i_pcie_usr_clk,                             // PCIE clock generated by end-point
    // PCIE EP - DMA engine interface
    input types_dma_pkg::dma64_in_type i_pcie_dmai,         // PCIE-EP to system DMA requests
    output types_dma_pkg::dma64_out_type o_pcie_dmao,       // System DMA responds to PCIE EP
    // DMA engine interface - System on Chip interface
    output types_pnp_pkg::dev_config_type o_xmst_cfg,       // PCIE DMA master interface descriptor
    input types_amba_pkg::axi4_master_in_type i_xmsti,
    output types_amba_pkg::axi4_master_out_type o_xmsto
);

import types_dma_pkg::*;
import types_pnp_pkg::*;
import types_amba_pkg::*;
import pcie_cfg_pkg::*;
import pcie_dma_pkg::*;

logic [TXFIFO_WIDTH-1:0] wb_txfifo_payload_i;
logic [TXFIFO_WIDTH-1:0] wb_txfifo_payload_o;
logic w_txfifo_full;
logic w_txfifo_empty;
logic w_txfifo_rd;
logic [RXFIFO_WIDTH-1:0] wb_rxfifo_payload_i;
logic [RXFIFO_WIDTH-1:0] wb_rxfifo_payload_o;
logic w_rxfifo_full;
logic w_rxfifo_empty;
logic w_rxfifo_wr;

// PCIE EP -> DMA
cdc_afifo #(
    .abits(CFG_PCIE_DMAFIFO_DEPTH),
    .dbits(TXFIFO_WIDTH)
) txfifo (
    .i_wclk(i_pcie_usr_clk),
    .i_wrstn(i_sys_nrst),
    .i_wr(i_pcie_dmai.tx_valid),
    .i_wdata(wb_txfifo_payload_i),
    .o_wfull(w_txfifo_full),
    .i_rclk(i_sys_clk),
    .i_rrstn(i_sys_nrst),
    .i_rd(w_txfifo_rd),
    .o_rdata(wb_txfifo_payload_o),
    .o_rempty(w_txfifo_empty)
);
// DMA -> PCIE EP
cdc_afifo #(
    .abits(CFG_PCIE_DMAFIFO_DEPTH),
    .dbits(RXFIFO_WIDTH)
) rxfifo (
    .i_wclk(i_pcie_usr_clk),
    .i_wrstn(i_sys_nrst),
    .i_wr(w_rxfifo_wr),
    .i_wdata(wb_rxfifo_payload_i),
    .o_wfull(w_rxfifo_full),
    .i_rclk(i_sys_clk),
    .i_rrstn(i_sys_nrst),
    .i_rd(i_pcie_dmai.rx_ready),
    .o_rdata(wb_rxfifo_payload_o),
    .o_rempty(w_rxfifo_empty)
);

always_comb
begin: comb_proc
    dev_config_type vb_xmst_cfg;
    logic [63:0] vb_tx_data;
    logic [7:0] vb_tx_strob;
    logic v_tx_last;
    logic [63:0] vb_rx_data;
    logic v_rx_last;

    vb_xmst_cfg = dev_config_none;
    vb_tx_data = 64'd0;
    vb_tx_strob = 8'd0;
    v_tx_last = 1'b0;
    vb_rx_data = 64'd0;
    v_rx_last = 1'b0;

    vb_xmst_cfg.descrsize = PNP_CFG_DEV_DESCR_BYTES;
    vb_xmst_cfg.descrtype = PNP_CFG_TYPE_MASTER;
    vb_xmst_cfg.vid = VENDOR_OPTIMITECH;
    vb_xmst_cfg.did = OPTIMITECH_PCIE_DMA;

    // TxFIFO inputs/outputs:
    wb_txfifo_payload_i = {i_pcie_dmai.tx_data,
            i_pcie_dmai.tx_strob,
            i_pcie_dmai.tx_last};

    vb_tx_data = wb_txfifo_payload_i[72: 9];
    vb_tx_strob = wb_txfifo_payload_i[8: 1];
    v_tx_last = wb_txfifo_payload_i[0];

    // RxFIFO inputs/outputs:
    wb_rxfifo_payload_i = {vb_rx_data,
            v_rx_last};

    o_pcie_dmao.rx_data = wb_rxfifo_payload_o[64: 1];
    o_pcie_dmao.rx_last = wb_rxfifo_payload_o[0];

    o_pcie_dmao.rx_valid = (~w_rxfifo_empty);
    o_pcie_dmao.tx_ready = (~w_txfifo_full);
    o_pcie_dmao.busy = 1'b0;
    w_txfifo_rd = 1'b1;
    o_xmst_cfg = vb_xmst_cfg;
    o_xmsto = axi4_master_out_none;
end: comb_proc

endmodule: pcie_dma
