// 
//  Copyright 2022 Sergey Khabarov, sergeykhbr@gmail.com
// 
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
// 

`timescale 1ps / 1ps

module pcie_app #(
  parameter logic async_reset = 1'b0,
  parameter C_DATA_WIDTH = 64,            // RX/TX interface data width

  // Do not override parameters below this line
  parameter KEEP_WIDTH = C_DATA_WIDTH / 8              // TSTRB width
) (
    input logic i_nrst,                                     // System Reset: active LOW
    input logic i_clk,                                      // System bus clock
    input logic i_pcie_phy_clk,                             // PCIE clock generated by end-point
    // PCIE EP - DMA engine interface
    input logic [15:0] i_pcie_completer_id,                 // Bus, Device, Function
    output logic [3:0] o_dma_state,                         // State machine debug output, connected to APB controller
    input types_dma_pkg::pcie_dma64_in_type i_pcie_dmai,    // PCIE-EP to system DMA requests
    output types_dma_pkg::pcie_dma64_out_type o_pcie_dmao,  // System DMA responds to PCIE EP
    // DMA engine interface - System on Chip interface
    output types_pnp_pkg::dev_config_type o_xmst_cfg,       // PCIE DMA master interface descriptor
    input types_amba_pkg::axi4_master_in_type i_xmsti,
    output types_amba_pkg::axi4_master_out_type o_xmsto,
    // Debug signals:
    output types_dma_pkg::pcie_dma64_in_type o_dbg_pcie_dmai
);

import types_dma_pkg::*;
import types_pnp_pkg::*;
import types_amba_pkg::*;
import pcie_cfg_pkg::*;
import pcie_dma_pkg::*;

  //----------------------------------------------------------------------------------------------------------------//
  // PCIe Block EP Tieoffs - Example PIO doesn't support the following inputs                                       //
  //----------------------------------------------------------------------------------------------------------------//

//  assign s_axis_tx_tuser[0] = 1'b0;                // Unused for V6
//  assign s_axis_tx_tuser[1] = 1'b0;                // Error forward packet
//  assign s_axis_tx_tuser[2] = 1'b0;                // Stream packet


//  wire [15:0] cfg_completer_id      = { i_cfg_bus_number, i_cfg_device_number, i_cfg_function_number };
//  wire  s_axis_tx_tready_i ;
//  assign s_axis_tx_tready_i = s_axis_tx_tready;
  wire [21:0] m_axis_rx_tuser;
  assign m_axis_rx_tuser = {'0, i_pcie_dmai.bar_hit, i_pcie_dmai.ecrc_err, i_pcie_dmai.err_fwd};

  assign o_xmst_cfg = dev_config_none;
  assign o_xmsto = axi4_master_out_none;
  assign o_dma_state = '0;
  assign o_dbg_pcie_dmai = pcie_dma64_in_none;


  //----------------------------------------------------------------------------------------------------------------//

  pcie_io  #(

    .C_DATA_WIDTH( C_DATA_WIDTH ),
    .KEEP_WIDTH( KEEP_WIDTH )

  ) PIO (

    .i_clk( i_clk ),
    .i_user_clk ( i_pcie_phy_clk ), //user_clk ),                         // I
    .i_user_reset ( ~i_nrst ), //user_reset ),                     // I
    .i_user_lnk_up ( i_nrst ), //i_user_lnk_up ),                   // I

    .i_s_axis_tx_tready ( i_pcie_dmai.ready ), //s_axis_tx_tready_i ),       // I
    .o_s_axis_tx_tdata  ( o_pcie_dmao.data ), //s_axis_tx_tdata ),          // O
    .o_s_axis_tx_tkeep  ( o_pcie_dmao.strob ), //s_axis_tx_tkeep ),          // O
    .o_s_axis_tx_tlast  ( o_pcie_dmao.last ), //s_axis_tx_tlast ),          // O
    .o_s_axis_tx_tvalid ( o_pcie_dmao.valid ), //s_axis_tx_tvalid ),         // O
    .o_tx_src_dsc       ( ), //s_axis_tx_tuser[3] ),       // O  unused assigned to 1'b0

    .i_m_axis_rx_tdata ( i_pcie_dmai.data ), //m_axis_rx_tdata ),           // I
    .i_m_axis_rx_tkeep ( i_pcie_dmai.strob ), //m_axis_rx_tkeep ),           // I
    .i_m_axis_rx_tlast ( i_pcie_dmai.last ), //m_axis_rx_tlast ),           // I
    .i_m_axis_rx_tvalid( i_pcie_dmai.valid ), //m_axis_rx_tvalid ),          // I
    .o_m_axis_rx_tready( o_pcie_dmao.ready ), //m_axis_rx_tready ),          // O
    .i_m_axis_rx_tuser ( m_axis_rx_tuser ),            // I

    .i_cfg_to_turnoff ( 1'b0 ), //i_cfg_to_turnoff ),             // I
    .o_cfg_turnoff_ok ( ),//o_cfg_turnoff_ok ),             // O
    .i_cfg_completer_id ( i_pcie_completer_id ) //cfg_completer_id ),         // I [15:0]
  );

endmodule // pcie_app
